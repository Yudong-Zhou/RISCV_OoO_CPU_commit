// module for Unified_Issue_Queue of Out-of-Order Processor
//
// Author: Yudong Zhou
//
// Create date: 11/9/2024
//
`timescale 1ns/1ps

module moduleName (
    ports
);
    
endmodule